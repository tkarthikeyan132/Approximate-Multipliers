

module AppHalfAdder(q0, p0, p1); 

input p0, p1;
output q0;

or or_1(q0, p0, p1);

endmodule
