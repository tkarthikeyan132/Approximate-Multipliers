

module Comp2p1(w0, p0, p1); // {p0+p1}

input p0, p1;
output w0;

or or_1(w0, p0, p1);

endmodule
